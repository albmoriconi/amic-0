--------------------------------------------------------------------------VHDL--
-- Copyright (C) 2019 Alberto Moriconi
--
-- This program is free software: you can redistribute it and/or modify it under
-- the terms of the GNU General Public License as published by the Free Software
-- Foundation, either version 3 of the License, or (at your option) any later
-- version.
--
-- This program is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS
-- FOR A PARTICULAR PURPOSE. See the GNU General Public License for more
-- details.
--
-- You should have received a copy of the GNU General Public License along with
-- this program. If not, see <http://www.gnu.org/licenses/>.
--------------------------------------------------------------------------------
--! @file control_store.vhd
--! @author Alberto Moriconi
--! @date 2019-05-11
--! @brief Processor control store
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.common_defs.all;

--! Processor control store

--! The control store is a ROM used to store the processor microprogram.
entity control_store is
  port (
    --! Address of the desired word
    address : in  ctrl_str_addr_type;
    --! Content of the addressed word
    word    : out ctrl_str_word_type;
    );
end entity control_store;

--! Dataflow architecture for the control store
architecture dataflow of control_store is

  -- Constants
  constant words : ctrl_str_type := (
--BEGIN_WORDS_ENTRY
    0      => "000000110111000000000000000000000000",
    1      => "010111100111000000000000000000000000",
    2      => "000000000000000000000000000000000000",
    3      => "000000000000000000000000000000000000",
    4      => "000000000000000000000000000000000000",
    5      => "000000000000000000000000000000000000",
    6      => "000000000100010000100000010101100001",
    7      => "000001000100000000100000010101100000",
    8      => "000001001100010000100000010101100000",
    9      => "000000110111000000000000000000000000",
    10     => "000000000000000000000000000000000000",
    11     => "000000000000000000000000000000000000",
    12     => "000000000000000000000000000000000000",
    13     => "000000000000000000000000000000000000",
    14     => "000000000000000000000000000000000000",
    15     => "000000000000000000000000000000000000",
    16     => "000010001001000010010000010101100000",
    17     => "000010010100010000100000010101100000",
    18     => "000000110010000101000010000101000000",
    19     => "000000000000000000000000000000000000",
    20     => "000000000000000000000000000000000000",
    21     => "000010110101000000000000100101000000",
    22     => "000010111110001010000000000111100000",
    23     => "000011000001000010010000010101100000",
    24     => "000011001100010100100000010101100000",
    25     => "000000110111000000000010000101000000",
    26     => "000000000000000000000000000000000000",
    27     => "000000000000000000000000000000000000",
    28     => "000000000000000000000000000000000000",
    29     => "000000000000000000000000000000000000",
    30     => "000000000000000000000000000000000000",
    31     => "000000000000000000000000000000000000",
    32     => "000100001100010000100000010101100000",
    33     => "000100010110000000000000100101001000",
    34     => "000100011110000000000000100111000000",
    35     => "000010111011001010000000000111100000",
    36     => "000000000000000000000000000000000000",
    37     => "000000000000000000000000000000000000",
    38     => "000000000000000000000000000000000000",
    39     => "000000000000000000000000000000000000",
    40     => "000000000000000000000000000000000000",
    41     => "000000000000000000000000000000000000",
    42     => "000000000000000000000000000000000000",
    43     => "000000000000000000000000000000000000",
    44     => "000000000000000000000000000000000000",
    45     => "000000000000000000000000000000000000",
    46     => "000000000000000000000000000000000000",
    47     => "000000000000000000000000000000000000",
    48     => "000000000000000000000000000000000000",
    49     => "000000000000000000000000000000000000",
    50     => "000000000000000000000000000000000000",
    51     => "000000000000000000000000000000000000",
    52     => "000000000000000000000000000000000000",
    53     => "000000000000000000000000000000000000",
    54     => "000110111101000000000000100101000000",
    55     => "000111000110000010000000000111100000",
    56     => "000111001111000101000000000101000000",
    57     => "000111010001001010010000001101100000",
    58     => "000111011100010000100000010101100000",
    59     => "000000110111000000000010000101000000",
    60     => "000000000000000000000000000000000000",
    61     => "000000000000000000000000000000000000",
    62     => "000000000000000000000000000000000000",
    63     => "000000000000000000000000000000000000",
    64     => "000000000000000000000000000000000000",
    65     => "000000000000000000000000000000000000",
    66     => "000000000000000000000000000000000000",
    67     => "000000000000000000000000000000000000",
    68     => "000000000000000000000000000000000000",
    69     => "000000000000000000000000000000000000",
    70     => "000000000000000000000000000000000000",
    71     => "000000000000000000000000000000000000",
    72     => "000000000000000000000000000000000000",
    73     => "000000000000000000000000000000000000",
    74     => "000000000000000000000000000000000000",
    75     => "000000000000000000000000000000000000",
    76     => "000000000000000000000000000000000000",
    77     => "000000000000000000000000000000000000",
    78     => "000000000000000000000000000000000000",
    79     => "000000000000000000000000000000000000",
    80     => "000000000000000000000000000000000000",
    81     => "000000000000000000000000000000000000",
    82     => "000000000000000000000000000000000000",
    83     => "000000000000000000000000000000000000",
    84     => "000000000000000000000000000000000000",
    85     => "000000000000000000000000000000000000",
    86     => "000000000000000000000000000000000000",
    87     => "001011000001000010010000010101100000",
    88     => "000000110111000101000000000101000000",
    89     => "001011010001001010010000001101100000",
    90     => "001011011111000000000000000000000000",
    91     => "000000110111000000000010000101000000",
    92     => "001011101001001010010000001101100000",
    93     => "001011110111000000000000100101000000",
    94     => "000000110111000101000010011111100000",
    95     => "001100000001001010000000001101100000",
    96     => "001100001001000010000000000101000000",
    97     => "001100010111000100000000100101000000",
    98     => "001100011111000001000000000101000000",
    99     => "001100100001000110000000001101100000",
    100    => "000000110111000000000010000011000000",
    101    => "001100110001001010010000001101100000",
    102    => "001100111111000000000000100101000000",
    103    => "000000110111000101000010000111100000",
    104    => "000000000000000000000000000000000000",
    105    => "000000000000000000000000000000000000",
    106    => "000000000000000000000000000000000000",
    107    => "000000000000000000000000000000000000",
    108    => "000000000000000000000000000000000000",
    109    => "000000000000000000000000000000000000",
    110    => "000000000000000000000000000000000000",
    111    => "000000000000000000000000000000000000",
    112    => "000000000000000000000000000000000000",
    113    => "000000000000000000000000000000000000",
    114    => "000000000000000000000000000000000000",
    115    => "000000000000000000000000000000000000",
    116    => "000000000000000000000000000000000000",
    117    => "000000000000000000000000000000000000",
    118    => "000000000000000000000000000000000000",
    119    => "000000000000000000000000000000000000",
    120    => "000000000000000000000000000000000000",
    121    => "000000000000000000000000000000000000",
    122    => "000000000000000000000000000000000000",
    123    => "000000000000000000000000000000000000",
    124    => "000000000000000000000000000000000000",
    125    => "000000000000000000000000000000000000",
    126    => "001111111001001010010000001101100000",
    127    => "010000000111000000000000100101000000",
    128    => "000000110111000101000010000110000000",
    129    => "000000000000000000000000000000000000",
    130    => "000000000000000000000000000000000000",
    131    => "000000000000000000000000000000000000",
    132    => "010000101101000000000000100101000000",
    133    => "010000110110001010000000000111100000",
    134    => "010000111100010000100000010101100000",
    135    => "010001000111000000000000100101000000",
    136    => "010001001100010000100000010101100000",
    137    => "000000110010000101000000000111100000",
    138    => "000000000000000000000000000000000000",
    139    => "000000000000000000000000000000000000",
    140    => "000000000000000000000000000000000000",
    141    => "000000000000000000000000000000000000",
    142    => "000000000000000000000000000000000000",
    143    => "000000000000000000000000000000000000",
    144    => "000000000000000000000000000000000000",
    145    => "000000000000000000000000000000000000",
    146    => "000000000000000000000000000000000000",
    147    => "000000000000000000000000000000000000",
    148    => "000000000000000000000000000000000000",
    149    => "000000000000000000000000000000000000",
    150    => "000000000000000000000000000000000000",
    151    => "000000000000000000000000000000000000",
    152    => "000000000000000000000000000000000000",
    153    => "010011010001001010010000001101100000",
    154    => "010011011111000000000001000101000000",
    155    => "010011100111000000000010000101000000",
    156    => "000000111000100000000000000101000100",
    157    => "010011110001001010010000001101100000",
    158    => "010011111111000000000001000101000000",
    159    => "010100000111000000000010000101000000",
    160    => "000000111000100000000000000101000010",
    161    => "010100010001001010010000001101100000",
    162    => "010100011001000010010000001101100000",
    163    => "010100100111001000000000100101000000",
    164    => "010100101111000000000001000101000000",
    165    => "010100110111000000000010000101000000",
    166    => "000000111000100000000000011111100100",
    167    => "010101000100000000000001001101100000",
    168    => "010101001100010000100000010101100000",
    169    => "010101010010000000000000100101001000",
    170    => "010101011110000000000000100111000000",
    171    => "010101100000110000100000000111100000",
    172    => "000000110111000000000000000000000000",
    173    => "010101110101001010010000000101000000",
    174    => "010101111111000000000000000000000000",
    175    => "010110000111001010001000000101000000",
    176    => "010110001101000010000000010101100000",
    177    => "010110010111011000100000000101000000",
    178    => "010110011001000010000000000101000000",
    179    => "010110100111000000001000000101000000",
    180    => "010110101111000101000000000101000000",
    181    => "000000110100000000000000001101100100",
    182    => "010110111001001010010000001101100000",
    183    => "010111000111000000000000100101000000",
    184    => "000000110111000101000010000111000000",
    185    => "010111010100010000100000010101100000",
    186    => "010111011110000000000000100101001000",
    187    => "010111100110000000000000100111000000",
    188    => "010111101011001010000000000111100000",
    189    => "010111110100000000000001010101100000",
    190    => "010111111111010000100000000101000000",
    191    => "011000000100010000100000010101100000",
    192    => "011000001110000000000000100101001000",
    193    => "011000010110000000000000100111000000",
    194    => "011000011100010000100000010101100000",
    195    => "011000100001000000000010011111100000",
    196    => "011000101111000010000010010101100000",
    197    => "011000110100010000100000010101100000",
    198    => "011000111110000000000000100101001000",
    199    => "011001000110000000000000100111000000",
    200    => "011001001001000101000000010111100000",
    201    => "011001010111000010010000000101000000",
    202    => "011001011000100101000000000101000000",
    203    => "011001100001000010010000010101100000",
    204    => "011001101101000101000000000101000000",
    205    => "011001110100010000100000010101100000",
    206    => "000000110111000000001000000101000000",
    207    => "100000000100010000100000010101100001",
    208    => "000000000000000000000000000000000000",
    209    => "000000000000000000000000000000000000",
    210    => "000000000000000000000000000000000000",
    211    => "000000000000000000000000000000000000",
    212    => "000000000000000000000000000000000000",
    213    => "000000000000000000000000000000000000",
    214    => "000000000000000000000000000000000000",
    215    => "000000000000000000000000000000000000",
    216    => "000000000000000000000000000000000000",
    217    => "000000000000000000000000000000000000",
    218    => "000000000000000000000000000000000000",
    219    => "000000000000000000000000000000000000",
    220    => "000000000000000000000000000000000000",
    221    => "000000000000000000000000000000000000",
    222    => "000000000000000000000000000000000000",
    223    => "000000000000000000000000000000000000",
    224    => "000000000000000000000000000000000000",
    225    => "000000000000000000000000000000000000",
    226    => "000000000000000000000000000000000000",
    227    => "000000000000000000000000000000000000",
    228    => "000000000000000000000000000000000000",
    229    => "000000000000000000000000000000000000",
    230    => "000000000000000000000000000000000000",
    231    => "000000000000000000000000000000000000",
    232    => "000000000000000000000000000000000000",
    233    => "000000000000000000000000000000000000",
    234    => "000000000000000000000000000000000000",
    235    => "000000000000000000000000000000000000",
    236    => "000000000000000000000000000000000000",
    237    => "000000000000000000000000000000000000",
    238    => "000000000000000000000000000000000000",
    239    => "000000000000000000000000000000000000",
    240    => "000000000000000000000000000000000000",
    241    => "000000000000000000000000000000000000",
    242    => "000000000000000000000000000000000000",
    243    => "000000000000000000000000000000000000",
    244    => "000000000000000000000000000000000000",
    245    => "000000000000000000000000000000000000",
    246    => "000000000000000000000000000000000000",
    247    => "000000000000000000000000000000000000",
    248    => "000000000000000000000000000000000000",
    249    => "000000000000000000000000000000000000",
    250    => "000000000000000000000000000000000000",
    251    => "000000000000000000000000000000000000",
    252    => "000000000000000000000000000000000000",
    253    => "000000000000000000000000000000000000",
    254    => "000000000000000000000000000000000000",
    255    => "000000000000000000000000000000000000",
    256    => "000000000000000000000000000000000000",
    257    => "000000000000000000000000000000000000",
    258    => "000000000000000000000000000000000000",
    259    => "000000000000000000000000000000000000",
    260    => "000000000000000000000000000000000000",
    261    => "000000000000000000000000000000000000",
    262    => "100000110111000000000000000000000000",
    263    => "010101000100010000000001001101100000",
    264    => "000000000000000000000000000000000000",
    265    => "000000000000000000000000000000000000",
    266    => "000000000000000000000000000000000000",
    267    => "000000000000000000000000000000000000",
    268    => "000000000000000000000000000000000000",
    269    => "000000000000000000000000000000000000",
    270    => "000000000000000000000000000000000000",
    271    => "000000000000000000000000000000000000",
    272    => "000000000000000000000000000000000000",
    273    => "000000000000000000000000000000000000",
    274    => "000000000000000000000000000000000000",
    275    => "000000000000000000000000000000000000",
    276    => "000000000000000000000000000000000000",
    277    => "100010110100010000100000010101100000",
    278    => "100010111110000000000000100101001000",
    279    => "100011000110000000000000100111000000",
    280    => "000010111101001010000000000111100000",
    281    => "000000000000000000000000000000000000",
    282    => "000000000000000000000000000000000000",
    283    => "000000000000000000000000000000000000",
    284    => "000000000000000000000000000000000000",
    285    => "000000000000000000000000000000000000",
    286    => "000000000000000000000000000000000000",
    287    => "000000000000000000000000000000000000",
    288    => "000000000000000000000000000000000000",
    289    => "000000000000000000000000000000000000",
    290    => "000000000000000000000000000000000000",
    291    => "000000000000000000000000000000000000",
    292    => "000000000000000000000000000000000000",
    293    => "000000000000000000000000000000000000",
    294    => "000000000000000000000000000000000000",
    295    => "000000000000000000000000000000000000",
    296    => "000000000000000000000000000000000000",
    297    => "000000000000000000000000000000000000",
    298    => "000000000000000000000000000000000000",
    299    => "000000000000000000000000000000000000",
    300    => "000000000000000000000000000000000000",
    301    => "000000000000000000000000000000000000",
    302    => "000000000000000000000000000000000000",
    303    => "000000000000000000000000000000000000",
    304    => "000000000000000000000000000000000000",
    305    => "000000000000000000000000000000000000",
    306    => "000000000000000000000000000000000000",
    307    => "000000000000000000000000000000000000",
    308    => "000000000000000000000000000000000000",
    309    => "000000000000000000000000000000000000",
    310    => "100110111100010000100000010101100000",
    311    => "100111000110000000000000100101001000",
    312    => "100111001110000000000000100111000000",
    313    => "000111000101000010000000000111100000",
    314    => "000000000000000000000000000000000000",
    315    => "000000000000000000000000000000000000",
    316    => "000000000000000000000000000000000000",
    317    => "000000000000000000000000000000000000",
    318    => "000000000000000000000000000000000000",
    319    => "000000000000000000000000000000000000",
    320    => "000000000000000000000000000000000000",
    321    => "000000000000000000000000000000000000",
    322    => "000000000000000000000000000000000000",
    323    => "000000000000000000000000000000000000",
    324    => "000000000000000000000000000000000000",
    325    => "000000000000000000000000000000000000",
    326    => "000000000000000000000000000000000000",
    327    => "000000000000000000000000000000000000",
    328    => "000000000000000000000000000000000000",
    329    => "000000000000000000000000000000000000",
    330    => "000000000000000000000000000000000000",
    331    => "000000000000000000000000000000000000",
    332    => "000000000000000000000000000000000000",
    333    => "000000000000000000000000000000000000",
    334    => "000000000000000000000000000000000000",
    335    => "000000000000000000000000000000000000",
    336    => "000000000000000000000000000000000000",
    337    => "000000000000000000000000000000000000",
    338    => "000000000000000000000000000000000000",
    339    => "000000000000000000000000000000000000",
    340    => "000000000000000000000000000000000000",
    341    => "000000000000000000000000000000000000",
    342    => "000000000000000000000000000000000000",
    343    => "000000000000000000000000000000000000",
    344    => "000000000000000000000000000000000000",
    345    => "000000000000000000000000000000000000",
    346    => "000000000000000000000000000000000000",
    347    => "000000000000000000000000000000000000",
    348    => "000000000000000000000000000000000000",
    349    => "000000000000000000000000000000000000",
    350    => "000000000000000000000000000000000000",
    351    => "000000000000000000000000000000000000",
    352    => "000000000000000000000000000000000000",
    353    => "000000000000000000000000000000000000",
    354    => "000000000000000000000000000000000000",
    355    => "000000000000000000000000000000000000",
    356    => "000000000000000000000000000000000000",
    357    => "000000000000000000000000000000000000",
    358    => "000000000000000000000000000000000000",
    359    => "000000000000000000000000000000000000",
    360    => "000000000000000000000000000000000000",
    361    => "000000000000000000000000000000000000",
    362    => "000000000000000000000000000000000000",
    363    => "000000000000000000000000000000000000",
    364    => "000000000000000000000000000000000000",
    365    => "000000000000000000000000000000000000",
    366    => "000000000000000000000000000000000000",
    367    => "000000000000000000000000000000000000",
    368    => "000000000000000000000000000000000000",
    369    => "000000000000000000000000000000000000",
    370    => "000000000000000000000000000000000000",
    371    => "000000000000000000000000000000000000",
    372    => "000000000000000000000000000000000000",
    373    => "000000000000000000000000000000000000",
    374    => "000000000000000000000000000000000000",
    375    => "000000000000000000000000000000000000",
    376    => "000000000000000000000000000000000000",
    377    => "000000000000000000000000000000000000",
    378    => "000000000000000000000000000000000000",
    379    => "000000000000000000000000000000000000",
    380    => "000000000000000000000000000000000000",
    381    => "000000000000000000000000000000000000",
    382    => "000000000000000000000000000000000000",
    383    => "000000000000000000000000000000000000",
    384    => "000000000000000000000000000000000000",
    385    => "000000000000000000000000000000000000",
    386    => "000000000000000000000000000000000000",
    387    => "000000000000000000000000000000000000",
    388    => "000000000000000000000000000000000000",
    389    => "000000000000000000000000000000000000",
    390    => "000000000000000000000000000000000000",
    391    => "000000000000000000000000000000000000",
    392    => "000000000000000000000000000000000000",
    393    => "000000000000000000000000000000000000",
    394    => "000000000000000000000000000000000000",
    395    => "000000000000000000000000000000000000",
    396    => "000000000000000000000000000000000000",
    397    => "000000000000000000000000000000000000",
    398    => "000000000000000000000000000000000000",
    399    => "000000000000000000000000000000000000",
    400    => "000000000000000000000000000000000000",
    401    => "000000000000000000000000000000000000",
    402    => "000000000000000000000000000000000000",
    403    => "000000000000000000000000000000000000",
    404    => "000000000000000000000000000000000000",
    405    => "000000000000000000000000000000000000",
    406    => "000000000000000000000000000000000000",
    407    => "000000000000000000000000000000000000",
    408    => "000000000000000000000000000000000000",
    409    => "000000000000000000000000000000000000",
    410    => "000000000000000000000000000000000000",
    411    => "000000000000000000000000000000000000",
    412    => "000000000000000000000000000000000000",
    413    => "000000000000000000000000000000000000",
    414    => "000000000000000000000000000000000000",
    415    => "000000000000000000000000000000000000",
    416    => "000000000000000000000000000000000000",
    417    => "000000000000000000000000000000000000",
    418    => "000000000000000000000000000000000000",
    419    => "000000000000000000000000000000000000",
    420    => "000000000000000000000000000000000000",
    421    => "000000000000000000000000000000000000",
    422    => "000000000000000000000000000000000000",
    423    => "000000000000000000000000000000000000",
    424    => "000000000000000000000000000000000000",
    425    => "000000000000000000000000000000000000",
    426    => "000000000000000000000000000000000000",
    427    => "000000000000000000000000000000000000",
    428    => "000000000000000000000000000000000000",
    429    => "000000000000000000000000000000000000",
    430    => "000000000000000000000000000000000000",
    431    => "000000000000000000000000000000000000",
    432    => "000000000000000000000000000000000000",
    433    => "000000000000000000000000000000000000",
    434    => "000000000000000000000000000000000000",
    435    => "000000000000000000000000000000000000",
    436    => "000000000000000000000000000000000000",
    437    => "000000000000000000000000000000000000",
    438    => "000000000000000000000000000000000000",
    439    => "000000000000000000000000000000000000",
    440    => "000000000000000000000000000000000000",
    441    => "000000000000000000000000000000000000",
    442    => "000000000000000000000000000000000000",
    443    => "000000000000000000000000000000000000",
    444    => "000000000000000000000000000000000000",
    445    => "000000000000000000000000000000000000",
    446    => "000000000000000000000000000000000000",
    447    => "000000000000000000000000000000000000",
    448    => "000000000000000000000000000000000000",
    449    => "000000000000000000000000000000000000",
    450    => "000000000000000000000000000000000000",
    451    => "000000000000000000000000000000000000",
    452    => "000000000000000000000000000000000000",
    453    => "000000000000000000000000000000000000",
    454    => "000000000000000000000000000000000000",
    455    => "000000000000000000000000000000000000",
    456    => "000000000000000000000000000000000000",
    457    => "000000000000000000000000000000000000",
    458    => "000000000000000000000000000000000000",
    459    => "000000000000000000000000000000000000",
    460    => "000000000000000000000000000000000000",
    461    => "000000000000000000000000000000000000",
    462    => "000000000000000000000000000000000000",
    463    => "000000000000000000000000000000000000",
    464    => "000000000000000000000000000000000000",
    465    => "000000000000000000000000000000000000",
    466    => "000000000000000000000000000000000000",
    467    => "000000000000000000000000000000000000",
    468    => "000000000000000000000000000000000000",
    469    => "000000000000000000000000000000000000",
    470    => "000000000000000000000000000000000000",
    471    => "000000000000000000000000000000000000",
    472    => "000000000000000000000000000000000000",
    473    => "000000000000000000000000000000000000",
    474    => "000000000000000000000000000000000000",
    475    => "000000000000000000000000000000000000",
    476    => "000000000000000000000000000000000000",
    477    => "000000000000000000000000000000000000",
    478    => "000000000000000000000000000000000000",
    479    => "000000000000000000000000000000000000",
    480    => "000000000000000000000000000000000000",
    481    => "000000000000000000000000000000000000",
    482    => "000000000000000000000000000000000000",
    483    => "000000000000000000000000000000000000",
    484    => "000000000000000000000000000000000000",
    485    => "000000000000000000000000000000000000",
    486    => "000000000000000000000000000000000000",
    487    => "000000000000000000000000000000000000",
    488    => "000000000000000000000000000000000000",
    489    => "000000000000000000000000000000000000",
    490    => "000000000000000000000000000000000000",
    491    => "000000000000000000000000000000000000",
    492    => "000000000000000000000000000000000000",
    493    => "000000000000000000000000000000000000",
    494    => "000000000000000000000000000000000000",
    495    => "000000000000000000000000000000000000",
    496    => "000000000000000000000000000000000000",
    497    => "000000000000000000000000000000000000",
    498    => "000000000000000000000000000000000000",
    499    => "000000000000000000000000000000000000",
    500    => "000000000000000000000000000000000000",
    501    => "000000000000000000000000000000000000",
    502    => "000000000000000000000000000000000000",
    503    => "000000000000000000000000000000000000",
    504    => "000000000000000000000000000000000000",
    505    => "000000000000000000000000000000000000",
    506    => "000000000000000000000000000000000000",
    507    => "000000000000000000000000000000000000",
    508    => "000000000000000000000000000000000000",
    509    => "000000000000000000000000000000000000",
    510    => "000000000000000000000000000000000000",
    511    => "000000000000000000000000000000000000",
    others => (others => '0')
--END_WORDS_ENTRY
    );

begin  -- architecture dataflow

  word <= words(to_integer(unsigned(address)));

end architecture dataflow;
